`ifndef LIBHDL_GLOBAL
`define LIBHDL_GLOBAL
`defaultnettype none
`endif