`ifndef LIBHDL_TIMESCALE
`define LIBHDL_TIMESCALE
`timescale 1 ns / 1 ps
`endif