`ifndef LIBHDL_GLOBAL
`define LIBHDL_GLOBAL
`default_nettype none
`endif
